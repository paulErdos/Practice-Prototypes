Life Stage Group|Total Water (L/d)|Carbohydrate (g/d)|Total Fiber (g/d)|Fat (g/d)|Linoleic Acid (g/d)|α-Linolenic Acid (g/d)|Protein (g/d)
Infants 0–6 mo   |0.7|60 |ND|31|4.4|0.5|9.1
Infants 6–12 mo  |0.8|95 |ND|30|4.6|0.5|11.0
Children 1–3 y   |1.3|130|19|ND|7  |0.7|13
Children 4–8 y   |1.7|130|25|ND|10 |0.9|19
Males 9–13 y     |2.4|130|31|ND|12 |1.2|34
Males 14–18 y    |3.3|130|38|ND|16 |1.6|52
Males 19–30 y    |3.7|130|38|ND|17 |1.6|56
Males 31–50 y    |3.7|130|38|ND|17 |1.6|56
Males 51–70 y    |3.7|130|30|ND|14 |1.6|56
Males > 70 y     |3.7|130|30|ND|14 |1.6|56
Females 9–13 y   |2.1|130|26|ND|10 |1.0|34
Females 14–18 y  |2.3|130|26|ND|11 |1.1|46
Females 19–30 y  |2.7|130|25|ND|12 |1.1|46
Females 31–50 y  |2.7|130|25|ND|12 |1.1|46
Females 51–70 y  |2.7|130|21|ND|11 |1.1|46
Females > 70 y   |2.7|130|21|ND|11 |1.1|46
Pregnancy 14–18 y|3.0|175|28|ND|13 |1.4|71
Pregnancy 19–30 y|3.0|175|28|ND|13 |1.4|71
Pregnancy 31–50 y|3.0|175|28|ND|13 |1.4|71
Lactation 14–18 y|3.8|210|29|ND|13 |1.3|71
Lactation 19–30 y|3.8|210|29|ND|13 |1.3|71
Lactation 31–50 y|3.8|210|29|ND|13 |1.3|71
#
# Source: https://www.ncbi.nlm.nih.gov/books/NBK56068/table/summarytables.t4/?report=objectonly