Life Stage Group|Vitamin A (μg/d)|Vitamin C (mg/d)|Vitamin D (μg/d)|Vitamin E (mg/d)|Vitamin K (μg/d)|Thiamin (mg/d)|Riboflavin (mg/d)|Niacin (mg/d)|Vitamin B6 (mg/d)|Folate (μg/d)f|Vitamin B12 (μg/d)|Pantothenic Acid (mg/d)|Biotin (μg/d)|Choline (mg/d)
Infants 0–6 mo|400|40|10|4|2.0|0.2|0.3|2|0.1|65|0.4|1.7|5|125
Infants 6–12 mo|500|50|10|5|2.5|0.3|0.4|4|0.3|80|0.5|1.8|6|150
Children 1–3 y|300|15|15|6|30|0.5|0.5|6|0.5|150|0.9|2|8|200
Children 4–8 y|400|25|15|7|55|0.6|0.6|8|0.6|200|1.2|3|12|250
Males 9–13 y|600|45|15|11|60|0.9|0.9|12|1.0|300|1.8|4|20|375
Males 14–18 y|900|75|15|15|75|1.2|1.3|16|1.3|400|2.4|5|25|550
Males 19–30 y|900|90|15|15|120|1.2|1.3|16|1.3|400|2.4|5|30|550
Males 31–50 y|900|90|15|15|120|1.2|1.3|16|1.3|400|2.4|5|30|550
Males 51–70 y|900|90|15|15|120|1.2|1.3|16|1.7|400|2.4|5|30|550
Males > 70 y|900|90|20|15|120|1.2|1.3|16|1.7|400|2.4|5|30|550
Females 9–13 y|600|45|15|11|60|0.9|0.9|12|1.0|300|1.8|4|20|375
Females 14–18 y|700|65|15|15|75|1.0|1.0|14|1.2|400i|2.4|5|25|400
Females 19–30 y|700|75|15|15|90|1.1|1.1|14|1.3|400i|2.4|5|30|425
Females 31–50 y|700|75|15|15|90|1.1|1.1|14|1.3|400i|2.4|5|30|425
Females 51–70 y|700|75|15|15|90|1.1|1.1|14|1.5|400|2.4|5|30|425
Females > 70 y|700|75|20|15|90|1.1|1.1|14|1.5|400|2.4|5|30|425
Pregnancy 14–18 y|750|80|15|15|75|1.4|1.4|18|1.9|600j|2.6|6|30|450
Pregnancy 19–30 y|770|85|15|15|90|1.4|1.4|18|1.9|600j|2.6|6|30|450
Pregnancy 31–50 y|770|85|15|15|90|1.4|1.4|18|1.9|600j|2.6|6|30|450
Lactation 14–18 y|1,200|115|15|19|75|1.4|1.6|17|2.0|500|2.8|7|35|550
Lactation 19–30 y|1,300|120|15|19|90|1.4|1.6|17|2.0|500|2.8|7|35|550
Lactation 31–50 y|1,300|120|15|19|90|1.4|1.6|17|2.0|500|2.8|7|35|550
#
# source: https://www.ncbi.nlm.nih.gov/books/NBK56068/table/summarytables.t2/?report=objectonly