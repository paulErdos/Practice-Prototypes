Life Stage Group|Calcium (mg/d)|Chromium (μg/d)|Copper (μg/d)|Fluoride (mg/d)|Iodine (μg/d)|Iron (mg/d)|Magnesium (mg/d)|Manganese (mg/d)|Molybdenum (μg/d)|Phosphorus (mg/d)|Selenium (μg/d)|Zinc (mg/d)|Potassium (mg/d)|Sodium (mg/d)|Chloride (g/d)
Infants 0–6 mo|200|0.2|200|0.01|110|0.27|30|0.003|2|100|15|2|400|110|0.18
Infants7–12 mo|260|5.5|220|0.5|130|11|75|0.6|3|275|20|3|860|370|0.57
Children 1–3 y|700|11|340|0.7|90|7|80|1.2|17|460|20|3|2,000|800|1.5
Children 4–8 y|1,000|15|440|1|90|10|130|1.5|22|500|30|5|2,300|1,000|1.9
Males 9–13 y  |1,300|25|700|2|120|8|240|1.9|34|1,250|40|8|2,500|1,200|2.3
Males 14–18 y|1,300|35|890|3|150|11|410|2.2|43|1,250|55|11|3,000|1,500|2.3
Males 19–30 y|1,000|35|900|4|150|8|400|2.3|45|700|55|11|3,400|1,500|2.3
Males 31–50 y|1,000|35|900|4|150|8|420|2.3|45|700|55|11|3,400|1,500|2.3
Males 51–70 y|1,000|30|900|4|150|8|420|2.3|45|700|55|11|3,400|1,500|2.0
Males > 70 y|1,200|30|900|4|150|8|420|2.3|45|700|55|11|3,400|1,500|1.8
Females 9–13 y|1,300|21|700|2|120|8|240|1.6|34|1,250|40|8|2,300|1,200|2.3
Females 14–18 y|1,300|24|890|3|150|15|360|1.6|43|1,250|55|9|2,300|1,500|2.3
Females 19–30 y|1,000|25|900|3|150|18|310|1.8|45|700|55|8|2,600|1,500|2.3
Females 31–50 y|1,000|25|900|3|150|18|320|1.8|45|700|55|8|2,600|1,500|2.3
Females 51–70 y|1,200|20|900|3|150|8|320|1.8|45|700|55|8|2,600|1,500|2.0
Females > 70 y|1,200|20|900|3|150|8|320|1.8|45|700|55|8|2,600|1,500|1.8
Pregnancy 14–18 y|1,300|29|1,000|3|220|27|400|2.0|50|1,250|60|12|2,600|1,500|2.3
Pregnancy 19–30 y|1,000|30|1,000|3|220|27|350|2.0|50|700|60|11|2,900|1,500|2.3
Pregnancy 31–50 y|1,000|30|1,000|3|220|27|360|2.0|50|700|60|11|2,900|1,500|2.3
Lactation 14–18 y|1,300|44|1,300|3|290|10|360|2.6|50|1,250|70|13|2,500|1,500|2.3
Lactation 19–30 y|1,000|45|1,300|3|290|9|310|2.6|50|700|70|12|2,800|1,500|2.3
Lactation 31–50 y|1,000|45|1,300|3|290|9|320|2.6|50|700|70|12|2,800|1,500|2.3
#
# source: https://ods.od.nih.gov/HealthInformation/nutrientrecommendations.aspx
# source: www.ncbi.nlm.nih.gov/books/NBK545442/table/appJ_tab3/?report=objectonly